module wide_main(
    input[64:0] wide_input,
    output[64:0] wide_output
);
    assign wide_output = wide_input;
endmodule
