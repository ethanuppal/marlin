module very_wide_main(
    input[199:0] very_wide_input,
    output[199:0] very_wide_output
);
    assign very_wide_output = very_wide_input;
endmodule
